magic
tech sky130A
timestamp 1598183786
<< metal1 >>
rect 690 795 720 825
rect 690 750 720 780
rect 705 735 720 750
<< end >>

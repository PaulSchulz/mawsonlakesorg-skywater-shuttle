magic
tech sky130A
timestamp 1598363904
<< metal1 >>
rect 1655 700 1690 705
rect 1650 695 1695 700
rect 1645 685 1700 695
rect 1645 680 1660 685
rect 1640 670 1660 680
rect 1685 670 1700 685
rect 1640 665 1665 670
rect 1645 660 1670 665
rect 1645 655 1675 660
rect 1645 650 1680 655
rect 1640 645 1685 650
rect 1635 640 1690 645
rect 1635 635 1655 640
rect 1670 635 1695 640
rect 1635 620 1650 635
rect 1675 630 1700 635
rect 1675 625 1705 630
rect 1675 620 1710 625
rect 1635 615 1655 620
rect 1670 615 1710 620
rect 1635 610 1710 615
rect 1640 605 1710 610
rect 1645 600 1680 605
rect 1695 600 1710 605
<< end >>

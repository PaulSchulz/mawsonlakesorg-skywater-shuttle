magic
tech sky130A
timestamp 1598181805
<< metal1 >>
rect 1245 170 1260 255
rect 1275 170 1290 255
rect 1245 160 1290 170
rect 1250 155 1285 160
rect 1255 150 1280 155
<< end >>

magic
tech sky130A
timestamp 1598356319
<< metal1 >>
rect 1200 750 1260 765
<< end >>

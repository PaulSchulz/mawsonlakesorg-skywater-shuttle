magic
tech sky130A
timestamp 1598355775
<< metal1 >>
rect 1155 800 1170 815
rect 1140 785 1185 800
rect 1155 770 1170 785
<< end >>

magic
tech sky130A
magscale 1 2
timestamp 1598753609
use font_41  font_41_0 libraries/sky130_ml_xx_hd/mag
timestamp 1598685393
transform 1 0 0 0 1 60
box 0 0 90 210
use font_a  font_a_0 ~/Documents/git/mawsonlakesorg-skywater-shuttle/magic/lib/font-sky130
timestamp 1598165416
transform 1 0 0 0 1 60
box 0 0 90 150
use font_b  font_b_0 ~/Documents/git/mawsonlakesorg-skywater-shuttle/magic/lib/font-sky130
timestamp 1598177753
transform 1 0 0 0 1 60
box 120 0 210 210
use font_3E  font_3E_0 libraries/sky130_ml_xx_hd/mag
timestamp 1598360501
transform 1 0 401 0 1 -1730
box -270 1530 -180 1680
use font_3C  font_3C_0 libraries/sky130_ml_xx_hd/mag
timestamp 1598360344
transform 1 0 391 0 1 -1734
box -390 1530 -300 1680
use font_c  font_c_0 ~/Documents/git/mawsonlakesorg-skywater-shuttle/magic/lib/font-sky130
timestamp 1598177753
transform 1 0 0 0 1 60
box 240 0 330 150
use font_d  font_d_0 ~/Documents/git/mawsonlakesorg-skywater-shuttle/magic/lib/font-sky130
timestamp 1598177753
transform 1 0 0 0 1 60
box 360 0 450 210
use font_3D  font_3D_0 libraries/sky130_ml_xx_hd/mag
timestamp 1598360266
transform 1 0 436 0 1 -1682
box -150 1530 -30 1620
use font_e  font_e_0 ~/Documents/git/mawsonlakesorg-skywater-shuttle/magic/lib/font-sky130
timestamp 1598165416
transform 1 0 0 0 1 60
box 480 0 570 150
use font_f  font_f_0 ~/Documents/git/mawsonlakesorg-skywater-shuttle/magic/lib/font-sky130
timestamp 1598177753
transform 1 0 0 0 1 60
box 600 0 690 210
use font_g  font_g_0 ~/Documents/git/mawsonlakesorg-skywater-shuttle/magic/lib/font-sky130
timestamp 1598165416
transform 1 0 0 0 1 60
box 720 -60 810 150
use font_h  font_h_0 ~/Documents/git/mawsonlakesorg-skywater-shuttle/magic/lib/font-sky130
timestamp 1598177753
transform 1 0 0 0 1 60
box 840 0 930 210
use font_i  font_i_0 ~/Documents/git/mawsonlakesorg-skywater-shuttle/magic/lib/font-sky130
timestamp 1598177753
transform 1 0 0 0 1 60
box 960 0 1020 210
use font_j  font_j_0 ~/Documents/git/mawsonlakesorg-skywater-shuttle/magic/lib/font-sky130
timestamp 1598177753
transform 1 0 0 0 1 60
box 1050 -60 1110 210
use font_k  font_k_0 ~/Documents/git/mawsonlakesorg-skywater-shuttle/magic/lib/font-sky130
timestamp 1598165416
transform 1 0 0 0 1 60
box 1140 0 1230 210
use font_l  font_l_0 ~/Documents/git/mawsonlakesorg-skywater-shuttle/magic/lib/font-sky130
timestamp 1598177753
transform 1 0 0 0 1 60
box 1260 0 1290 210
use font_m  font_m_0 ~/Documents/git/mawsonlakesorg-skywater-shuttle/magic/lib/font-sky130
timestamp 1598177753
transform 1 0 0 0 1 60
box 1320 0 1470 150
use font_o  font_o_0 ~/Documents/git/mawsonlakesorg-skywater-shuttle/magic/lib/font-sky130
timestamp 1598165416
transform 1 0 0 0 1 60
box 1620 0 1710 150
use font_n  font_n_0 ~/Documents/git/mawsonlakesorg-skywater-shuttle/magic/lib/font-sky130
timestamp 1598165416
transform 1 0 0 0 1 60
box 1500 0 1590 150
use font_q  font_q_0 ~/Documents/git/mawsonlakesorg-skywater-shuttle/magic/lib/font-sky130
timestamp 1598177753
transform 1 0 0 0 1 60
box 1860 -60 1950 150
use font_p  font_p_0 ~/Documents/git/mawsonlakesorg-skywater-shuttle/magic/lib/font-sky130
timestamp 1598177753
transform 1 0 0 0 1 60
box 1740 -60 1830 150
use font_s  font_s_0 ~/Documents/git/mawsonlakesorg-skywater-shuttle/magic/lib/font-sky130
timestamp 1598165416
transform 1 0 0 0 1 60
box 2100 0 2190 150
use font_r  font_r_0 ~/Documents/git/mawsonlakesorg-skywater-shuttle/magic/lib/font-sky130
timestamp 1598165416
transform 1 0 0 0 1 60
box 1980 0 2070 150
use font_t  font_t_0 ~/Documents/git/mawsonlakesorg-skywater-shuttle/magic/lib/font-sky130
timestamp 1598177753
transform 1 0 0 0 1 60
box 2220 0 2310 180
use font_u  font_u_0 ~/Documents/git/mawsonlakesorg-skywater-shuttle/magic/lib/font-sky130
timestamp 1598177753
transform 1 0 0 0 1 60
box 2340 0 2430 150
use font_v  font_v_0 ~/Documents/git/mawsonlakesorg-skywater-shuttle/magic/lib/font-sky130
timestamp 1598177753
transform 1 0 0 0 1 60
box 2460 0 2550 150
use font_w  font_w_0 ~/Documents/git/mawsonlakesorg-skywater-shuttle/magic/lib/font-sky130
timestamp 1598166646
transform 1 0 0 0 1 60
box 2580 0 2730 150
use font_x  font_x_0 ~/Documents/git/mawsonlakesorg-skywater-shuttle/magic/lib/font-sky130
timestamp 1598177753
transform 1 0 0 0 1 60
box 2760 0 2850 150
use font_y  font_y_0 ~/Documents/git/mawsonlakesorg-skywater-shuttle/magic/lib/font-sky130
timestamp 1598177753
transform 1 0 0 0 1 60
box 2880 -60 2970 150
use font_z  font_z_0 ~/Documents/git/mawsonlakesorg-skywater-shuttle/magic/lib/font-sky130
timestamp 1598177753
transform 1 0 0 0 1 60
box 3000 0 3090 150
use font_24  font_24_0 libraries/sky130_ml_xx_hd/mag
timestamp 1598362656
transform 1 0 0 0 1 -840
box 3120 870 3210 1080
use font_2C  font_2C_0 libraries/sky130_ml_xx_hd/mag
timestamp 1598363612
transform 1 0 0 0 1 -840
box 3240 870 3300 960
use font_01F600  font_01F600_0 libraries/sky130_ml_xx_hd/mag
timestamp 1598364576
transform 1 0 0 0 1 -840
box 3330 900 3540 1070
use font_B  font_B_0 ~/Documents/git/mawsonlakesorg-skywater-shuttle/magic/lib/font-sky130
timestamp 1598181805
transform 1 0 0 0 1 60
box 120 300 210 510
use font_C  font_C_0 ~/Documents/git/mawsonlakesorg-skywater-shuttle/magic/lib/font-sky130
timestamp 1598181805
transform 1 0 0 0 1 60
box 240 300 330 510
use font_D  font_D_0 ~/Documents/git/mawsonlakesorg-skywater-shuttle/magic/lib/font-sky130
timestamp 1598181805
transform 1 0 120 0 1 60
box 240 300 330 510
use font_E  font_E_0 ~/Documents/git/mawsonlakesorg-skywater-shuttle/magic/lib/font-sky130
timestamp 1598181805
transform 1 0 0 0 1 60
box 480 300 570 510
use font_F  font_F_0 ~/Documents/git/mawsonlakesorg-skywater-shuttle/magic/lib/font-sky130
timestamp 1598181805
transform 1 0 0 0 1 60
box 600 300 690 510
use font_G  font_G_0 ~/Documents/git/mawsonlakesorg-skywater-shuttle/magic/lib/font-sky130
timestamp 1598181805
transform 1 0 0 0 1 60
box 720 300 810 510
use font_H  font_H_0 ~/Documents/git/mawsonlakesorg-skywater-shuttle/magic/lib/font-sky130
timestamp 1598181805
transform 1 0 0 0 1 60
box 840 300 930 510
use font_I  font_I_0 ~/Documents/git/mawsonlakesorg-skywater-shuttle/magic/lib/font-sky130
timestamp 1598181805
transform 1 0 0 0 1 60
box 960 300 1050 510
use font_K  font_K_0 ~/Documents/git/mawsonlakesorg-skywater-shuttle/magic/lib/font-sky130
timestamp 1598181805
transform 1 0 0 0 1 60
box 1200 300 1290 510
use font_J  font_J_0 ~/Documents/git/mawsonlakesorg-skywater-shuttle/magic/lib/font-sky130
timestamp 1598181805
transform 1 0 0 0 1 60
box 1080 300 1170 510
use font_L  font_L_0 ~/Documents/git/mawsonlakesorg-skywater-shuttle/magic/lib/font-sky130
timestamp 1598165416
transform 1 0 0 0 1 60
box 1320 300 1410 510
use font_M  font_M_0 ~/Documents/git/mawsonlakesorg-skywater-shuttle/magic/lib/font-sky130
timestamp 1598165416
transform 1 0 0 0 1 60
box 1440 300 1590 510
use font_A9  font_A9_0 libraries/sky130_ml_xx_hd/mag
timestamp 1598433283
transform 1 0 -240 0 1 -840
box 1710 1440 1920 1710
use font_N  font_N_0 ~/Documents/git/mawsonlakesorg-skywater-shuttle/magic/lib/font-sky130
timestamp 1598181805
transform 1 0 0 0 1 60
box 1620 300 1740 510
use font_P  font_P_0 ~/Documents/git/mawsonlakesorg-skywater-shuttle/magic/lib/font-sky130
timestamp 1598181805
transform 1 0 0 0 1 60
box 1890 300 1980 510
use font_O  font_O_0 ~/Documents/git/mawsonlakesorg-skywater-shuttle/magic/lib/font-sky130
timestamp 1598165416
transform 1 0 0 0 1 60
box 1770 300 1860 510
use font_40  font_at_0 libraries/sky130_ml_xx_hd/mag
timestamp 1598185717
transform 1 0 0 0 1 -840
box 1710 1440 1920 1710
use font_Q  font_Q_0 ~/Documents/git/mawsonlakesorg-skywater-shuttle/magic/lib/font-sky130
timestamp 1598181805
transform 1 0 0 0 1 60
box 2010 300 2100 510
use font_R  font_R_0 ~/Documents/git/mawsonlakesorg-skywater-shuttle/magic/lib/font-sky130
timestamp 1598181805
transform 1 0 0 0 1 60
box 2130 300 2220 510
use font_S  font_S_0 ~/Documents/git/mawsonlakesorg-skywater-shuttle/magic/lib/font-sky130
timestamp 1598181805
transform 1 0 0 0 1 60
box 2250 300 2340 510
use font_U  font_U_0 ~/Documents/git/mawsonlakesorg-skywater-shuttle/magic/lib/font-sky130
timestamp 1598181805
transform 1 0 0 0 1 60
box 2490 300 2580 510
use font_T  font_T_0 ~/Documents/git/mawsonlakesorg-skywater-shuttle/magic/lib/font-sky130
timestamp 1598181805
transform 1 0 0 0 1 60
box 2370 300 2460 510
use font_V  font_V_0 ~/Documents/git/mawsonlakesorg-skywater-shuttle/magic/lib/font-sky130
timestamp 1598181805
transform 1 0 0 0 1 60
box 2610 300 2700 510
use font_W  font_W_0 ~/Documents/git/mawsonlakesorg-skywater-shuttle/magic/lib/font-sky130
timestamp 1598181805
transform 1 0 0 0 1 60
box 2730 300 2880 510
use font_X  font_X_0 ~/Documents/git/mawsonlakesorg-skywater-shuttle/magic/lib/font-sky130
timestamp 1598181805
transform 1 0 0 0 1 60
box 2910 300 3000 510
use font_Y  font_Y_0 ~/Documents/git/mawsonlakesorg-skywater-shuttle/magic/lib/font-sky130
timestamp 1598181805
transform 1 0 0 0 1 60
box 3030 300 3120 510
use font_Z  font_Z_0 ~/Documents/git/mawsonlakesorg-skywater-shuttle/magic/lib/font-sky130
timestamp 1598181805
transform 1 0 0 0 1 60
box 3150 300 3240 510
use font_26  font_26_0 libraries/sky130_ml_xx_hd/mag
timestamp 1598363904
transform 1 0 0 0 1 -840
box 3270 1200 3420 1410
use font_3F  font_3F_0 libraries/sky130_ml_xx_hd/mag
timestamp 1598364457
transform 1 0 0 0 1 -840
box 3450 1200 3540 1410
use font_2E  font_2E_0 libraries/sky130_ml_xx_hd/mag
timestamp 1598165416
transform 1 0 -1920 0 1 660
box 3120 0 3180 60
use font_27  font_27_0 libraries/sky130_ml_xx_hd/mag
timestamp 1598355651
transform 1 0 0 0 1 -840
box 2040 1620 2100 1710
use font_21  font_21_0 libraries/sky130_ml_xx_hd/mag
timestamp 1598361454
transform 1 0 0 0 1 -840
box 1950 1500 2010 1710
use font_2D  font_2D_0 libraries/sky130_ml_xx_hd/mag
timestamp 1598355651
transform 1 0 0 0 1 -820
box 2130 1570 2250 1600
use font_2B  font_2B_0 libraries/sky130_ml_xx_hd/mag
timestamp 1598355775
transform 1 0 0 0 1 -820
box 2280 1540 2370 1630
use font_5F  font_5F_0 libraries/sky130_ml_xx_hd/mag
timestamp 1598356319
transform 1 0 0 0 1 -840
box 2400 1500 2520 1530
use font_5B  font_5B_0 libraries/sky130_ml_xx_hd/mag
timestamp 1598356361
transform 1 0 -120 0 1 -840
box 2670 1500 2760 1710
use font_5D  font_5D_0 libraries/sky130_ml_xx_hd/mag
timestamp 1598356419
transform 1 0 -120 0 1 -840
box 2790 1500 2880 1710
use font_5E  font_5E_0 libraries/sky130_ml_xx_hd/mag
timestamp 1598356481
transform 1 0 -120 0 1 -840
box 2910 1650 3000 1710
use font_23  font_23_0 libraries/sky130_ml_xx_hd/mag
timestamp 1598356557
transform 1 0 -120 0 1 -840
box 3030 1500 3180 1710
use font_60  font_60_0 libraries/sky130_ml_xx_hd/mag
timestamp 1598356612
transform 1 0 -120 0 1 -840
box 3210 1620 3270 1710
use font_2F  font_2F_0 libraries/sky130_ml_xx_hd/mag
timestamp 1598356782
transform 1 0 -120 0 1 -840
box 3300 1500 3390 1710
use font_25  font_25_0 libraries/sky130_ml_xx_hd/mag
timestamp 1598356858
transform 1 0 -120 0 1 -840
box 3420 1500 3570 1710
use font_7C  font_7C_0 libraries/sky130_ml_xx_hd/mag
timestamp 1598356911
transform 1 0 -120 0 1 -840
box 3600 1500 3630 1710
use font_7B  font_7B_0 libraries/sky130_ml_xx_hd/mag
timestamp 1598356953
transform 1 0 -120 0 1 -840
box 3660 1500 3750 1710
use font_7D  font_7D_0 libraries/sky130_ml_xx_hd/mag
timestamp 1598359058
transform 1 0 -120 0 1 -840
box 3780 1500 3870 1710
use font_7E  font_7E_0 libraries/sky130_ml_xx_hd/mag
timestamp 1598359164
transform 1 0 -120 0 1 -830
box 3900 1630 4050 1700
use font_22  font_22_0 libraries/sky130_ml_xx_hd/mag
timestamp 1598359472
transform -1 0 8130 0 1 -830
box 4080 1580 4170 1700
use font_2A  font_2A_0 libraries/sky130_ml_xx_hd/mag
timestamp 1598362535
transform 1 0 -10 0 1 -840
box 4090 1540 4220 1670
<< properties >>
string FIXED_BBOX -14 -854 104 -616
<< end >>

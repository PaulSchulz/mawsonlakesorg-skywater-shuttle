magic
tech sky130A
timestamp 1598165416
<< metal1 >>
rect 660 165 675 255
rect 660 150 705 165
<< end >>

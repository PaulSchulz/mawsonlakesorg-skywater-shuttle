magic
tech sky130A
timestamp 1598177753
<< metal1 >>
rect 1170 20 1185 75
rect 1200 20 1215 75
rect 1170 10 1215 20
rect 1175 5 1215 10
rect 1180 0 1215 5
<< end >>

magic
tech sky130A
timestamp 1598361454
<< metal1 >>
rect 975 795 1005 855
rect 975 750 1005 780
<< end >>

magic
tech sky130A
timestamp 1598177753
<< metal1 >>
rect 130 70 155 75
rect 125 65 160 70
rect 120 55 165 65
rect 120 20 135 55
rect 150 45 165 55
rect 150 20 165 25
rect 120 10 165 20
rect 125 5 160 10
rect 130 0 155 5
<< end >>

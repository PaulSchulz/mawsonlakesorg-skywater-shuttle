magic
tech sky130A
timestamp 1598356782
<< metal1 >>
rect 1680 840 1695 855
rect 1675 825 1695 840
rect 1670 820 1695 825
rect 1670 815 1690 820
rect 1665 810 1690 815
rect 1665 805 1685 810
rect 1660 800 1685 805
rect 1660 795 1680 800
rect 1655 790 1680 795
rect 1655 785 1675 790
rect 1650 780 1675 785
rect 1650 765 1670 780
rect 1650 750 1665 765
<< end >>

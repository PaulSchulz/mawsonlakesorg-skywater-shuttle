magic
tech sky130A
timestamp 1598362656
<< metal1 >>
rect 1575 525 1590 540
rect 1570 520 1605 525
rect 1565 515 1605 520
rect 1560 510 1605 515
rect 1560 495 1580 510
rect 1560 490 1595 495
rect 1565 485 1600 490
rect 1570 480 1605 485
rect 1585 465 1605 480
rect 1560 460 1605 465
rect 1560 455 1600 460
rect 1560 450 1595 455
rect 1575 435 1590 450
<< end >>

magic
tech sky130A
timestamp 1598181805
<< metal1 >>
rect 1575 240 1620 255
rect 1605 220 1620 240
rect 1600 215 1620 220
rect 1595 210 1620 215
rect 1590 205 1615 210
rect 1585 200 1610 205
rect 1580 195 1605 200
rect 1575 190 1600 195
rect 1575 185 1595 190
rect 1575 165 1590 185
rect 1575 150 1620 165
<< end >>

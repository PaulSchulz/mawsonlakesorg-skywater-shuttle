magic
tech sky130A
timestamp 1598181805
<< metal1 >>
rect 600 230 615 255
rect 630 230 645 255
rect 600 220 645 230
rect 600 210 640 220
rect 600 195 635 210
rect 600 185 640 195
rect 600 175 645 185
rect 600 150 615 175
rect 630 150 645 175
<< end >>

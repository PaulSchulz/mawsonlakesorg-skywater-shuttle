magic
tech sky130A
timestamp 1598165416
<< metal1 >>
rect 720 240 735 255
rect 780 240 795 255
rect 720 225 750 240
rect 765 225 795 240
rect 720 210 795 225
rect 720 150 735 210
rect 750 195 765 210
rect 780 150 795 210
<< end >>

magic
tech sky130A
timestamp 1598360344
<< metal1 >>
rect -165 835 -150 840
rect -170 830 -150 835
rect -175 825 -150 830
rect -180 820 -155 825
rect -185 815 -160 820
rect -190 810 -165 815
rect -195 795 -170 810
rect -190 790 -165 795
rect -185 785 -160 790
rect -180 780 -155 785
rect -175 775 -150 780
rect -170 770 -150 775
rect -165 765 -150 770
<< end >>

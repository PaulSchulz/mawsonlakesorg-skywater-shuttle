magic
tech sky130A
timestamp 1598359058
<< metal1 >>
rect 1890 850 1910 855
rect 1890 845 1915 850
rect 1890 835 1920 845
rect 1905 820 1920 835
rect 1905 810 1925 820
rect 1910 795 1935 810
rect 1905 785 1925 795
rect 1905 770 1920 785
rect 1890 760 1920 770
rect 1890 755 1915 760
rect 1890 750 1910 755
<< end >>

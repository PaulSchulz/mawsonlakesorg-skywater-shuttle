magic
tech sky130A
timestamp 1598177753
<< metal1 >>
rect 210 75 225 105
rect 190 70 225 75
rect 185 65 225 70
rect 180 55 225 65
rect 180 20 195 55
rect 210 20 225 55
rect 180 10 225 20
rect 185 5 225 10
rect 190 0 225 5
<< end >>

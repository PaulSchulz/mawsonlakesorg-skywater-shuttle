magic
tech sky130A
timestamp 1598181805
<< metal1 >>
rect 945 250 980 255
rect 945 245 985 250
rect 945 235 990 245
rect 945 200 960 235
rect 975 200 990 235
rect 945 190 990 200
rect 945 185 985 190
rect 945 180 980 185
rect 945 150 960 180
<< end >>

magic
tech sky130A
timestamp 1598359472
<< metal1 >>
rect 2040 790 2055 850
rect 2070 790 2085 850
<< end >>

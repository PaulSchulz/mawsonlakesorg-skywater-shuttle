magic
tech sky130A
timestamp 1598181805
<< metal1 >>
rect 1185 240 1230 255
rect 1200 150 1215 240
<< end >>

magic
tech sky130A
timestamp 1598361454
<< metal1 >>
rect 1570 550 1590 555
rect 1565 545 1590 550
rect 1560 535 1590 545
rect 1560 470 1575 535
rect 1560 460 1590 470
rect 1565 455 1590 460
rect 1570 450 1590 455
<< end >>

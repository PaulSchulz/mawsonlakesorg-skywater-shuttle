magic
tech sky130A
timestamp 1598182001
<< metal1 >>
rect 420 390 465 405
rect 450 300 465 390
<< end >>

magic
tech sky130A
timestamp 1598182001
<< metal1 >>
rect 360 390 405 405
rect 360 375 375 390
rect 360 360 405 375
rect 360 315 375 360
rect 390 315 405 360
rect 360 300 405 315
<< end >>

magic
tech sky130A
timestamp 1598182001
<< metal1 >>
rect 120 390 165 405
rect 150 375 165 390
rect 120 360 165 375
rect 120 315 135 360
rect 120 300 165 315
<< end >>

magic
tech sky130A
timestamp 1598361454
<< metal1 >>
rect 1605 550 1625 555
rect 1605 545 1630 550
rect 1605 535 1635 545
rect 1620 470 1635 535
rect 1605 460 1635 470
rect 1605 455 1630 460
rect 1605 450 1625 455
<< end >>

magic
tech sky130A
timestamp 1598356557
<< metal1 >>
rect 1530 825 1545 855
rect 1560 825 1575 855
rect 1515 810 1590 825
rect 1530 795 1545 810
rect 1560 795 1575 810
rect 1515 780 1590 795
rect 1530 750 1545 780
rect 1560 750 1575 780
<< end >>

magic
tech sky130A
timestamp 1598165416
<< metal1 >>
rect 1060 70 1095 75
rect 1055 65 1095 70
rect 1050 60 1095 65
rect 1050 45 1070 60
rect 1050 40 1085 45
rect 1055 35 1090 40
rect 1060 30 1095 35
rect 1075 15 1095 30
rect 1050 10 1095 15
rect 1050 5 1090 10
rect 1050 0 1085 5
<< end >>

magic
tech sky130A
timestamp 1598360501
<< metal1 >>
rect -135 835 -120 840
rect -135 830 -115 835
rect -135 825 -110 830
rect -130 820 -105 825
rect -125 815 -100 820
rect -120 810 -95 815
rect -115 795 -90 810
rect -120 790 -95 795
rect -125 785 -100 790
rect -130 780 -105 785
rect -135 775 -110 780
rect -135 770 -115 775
rect -135 765 -120 770
<< end >>

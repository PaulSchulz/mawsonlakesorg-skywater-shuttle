magic
tech sky130A
timestamp 1598685393
<< metal5 >>
rect -1495 98565 98705 98765
rect -1495 -1235 -1295 98565
rect 98505 -1235 98705 98565
rect -1495 -1435 98705 -1235
use font-sky130  font-sky130_0 ~/Documents/git/mawsonlakesorg-skywater-shuttle/magic
timestamp 1598532849
transform 1 0 0 0 1 -600
box -195 420 2105 855
use open-source-hardware  open-source-hardware_0
timestamp 1597969098
transform 1 0 -1195 0 1 -1030
box 0 -105 615 555
<< end >>

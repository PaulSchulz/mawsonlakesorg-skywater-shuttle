magic
tech sky130A
timestamp 1598177753
<< metal1 >>
rect 1500 60 1545 75
rect 1520 45 1545 60
rect 1515 40 1540 45
rect 1510 35 1535 40
rect 1505 30 1530 35
rect 1500 15 1525 30
rect 1500 0 1545 15
<< end >>

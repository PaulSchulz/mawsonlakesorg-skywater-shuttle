magic
tech sky130A
timestamp 1598356481
<< metal1 >>
rect 1470 840 1485 855
rect 1455 825 1500 840
<< end >>

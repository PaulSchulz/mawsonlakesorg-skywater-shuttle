magic
tech sky130A
timestamp 1598181805
<< metal1 >>
rect 370 250 395 255
rect 365 245 400 250
rect 360 235 405 245
rect 360 170 375 235
rect 390 225 405 235
rect 390 170 405 210
rect 360 160 405 170
rect 365 155 405 160
rect 370 150 405 155
<< end >>

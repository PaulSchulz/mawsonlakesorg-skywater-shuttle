magic
tech sky130A
timestamp 1597975676
<< metal1 >>
rect 255 540 330 555
rect 120 495 165 510
rect 105 480 195 495
rect 240 480 345 540
rect 420 495 465 510
rect 390 480 480 495
rect 105 465 210 480
rect 225 465 360 480
rect 375 465 480 480
rect 105 450 480 465
rect 120 420 465 450
rect 135 405 450 420
rect 150 390 440 405
rect 135 375 255 390
rect 330 375 450 390
rect 75 360 240 375
rect 345 360 510 375
rect 45 285 225 360
rect 360 285 525 360
rect 75 270 240 285
rect 345 270 510 285
rect 135 255 255 270
rect 150 240 255 255
rect 330 255 450 270
rect 330 240 435 255
rect 135 225 240 240
rect 120 210 240 225
rect 345 225 450 240
rect 345 210 465 225
rect 120 195 225 210
rect 105 180 225 195
rect 360 195 465 210
rect 360 180 480 195
rect 105 165 210 180
rect 375 165 480 180
rect 105 150 195 165
rect 390 150 480 165
rect 120 135 165 150
rect 420 135 465 150
rect 10 70 35 75
rect 70 70 95 75
rect 125 70 160 75
rect 180 70 215 75
rect 280 70 315 75
rect 340 70 365 75
rect 5 65 40 70
rect 65 65 100 70
rect 0 55 45 65
rect 0 20 15 55
rect 30 20 45 55
rect 0 10 45 20
rect 60 55 105 65
rect 60 20 75 55
rect 90 20 105 55
rect 60 10 105 20
rect 120 60 165 70
rect 120 45 135 60
rect 150 45 165 60
rect 120 35 165 45
rect 180 65 220 70
rect 275 65 315 70
rect 335 65 370 70
rect 180 55 225 65
rect 120 30 160 35
rect 120 15 135 30
rect 5 5 40 10
rect 60 5 100 10
rect 120 5 165 15
rect 10 0 35 5
rect 60 0 95 5
rect 125 0 165 5
rect 180 0 195 55
rect 210 0 225 55
rect 270 60 315 65
rect 270 45 290 60
rect 330 55 375 65
rect 270 40 305 45
rect 275 35 310 40
rect 280 30 315 35
rect 295 15 315 30
rect 270 10 315 15
rect 330 20 345 55
rect 360 20 375 55
rect 330 10 375 20
rect 390 20 405 75
rect 420 20 435 75
rect 390 10 435 20
rect 450 70 485 75
rect 520 70 545 75
rect 575 70 610 75
rect 450 65 490 70
rect 515 65 550 70
rect 450 55 495 65
rect 270 5 310 10
rect 335 5 370 10
rect 395 5 430 10
rect 270 0 305 5
rect 340 0 365 5
rect 400 0 425 5
rect 450 0 465 55
rect 480 45 495 55
rect 510 55 555 65
rect 510 20 525 55
rect 540 45 555 55
rect 570 60 615 70
rect 570 45 585 60
rect 600 45 615 60
rect 570 35 615 45
rect 570 30 610 35
rect 540 20 555 30
rect 510 10 555 20
rect 570 15 585 30
rect 515 5 550 10
rect 570 5 615 15
rect 520 0 545 5
rect 575 0 615 5
rect 60 -30 75 0
rect 270 -30 285 0
rect 60 -35 95 -30
rect 120 -35 160 -30
rect 180 -35 215 -30
rect 250 -35 285 -30
rect 60 -40 100 -35
rect 60 -50 105 -40
rect 120 -45 165 -35
rect 60 -105 75 -50
rect 90 -105 105 -50
rect 150 -60 165 -45
rect 120 -75 165 -60
rect 120 -90 135 -75
rect 150 -90 165 -75
rect 120 -100 165 -90
rect 125 -105 165 -100
rect 180 -40 220 -35
rect 245 -40 285 -35
rect 180 -50 225 -40
rect 180 -105 195 -50
rect 210 -60 225 -50
rect 240 -50 285 -40
rect 240 -85 255 -50
rect 270 -85 285 -50
rect 240 -95 285 -85
rect 300 -85 315 -30
rect 330 -85 345 -30
rect 360 -85 375 -30
rect 390 -35 430 -30
rect 450 -35 485 -30
rect 515 -35 550 -30
rect 390 -45 435 -35
rect 420 -60 435 -45
rect 395 -65 435 -60
rect 300 -95 375 -85
rect 390 -75 435 -65
rect 390 -90 405 -75
rect 420 -90 435 -75
rect 245 -100 285 -95
rect 305 -100 370 -95
rect 390 -100 435 -90
rect 250 -105 285 -100
rect 310 -105 330 -100
rect 345 -105 365 -100
rect 395 -105 435 -100
rect 450 -40 490 -35
rect 450 -50 495 -40
rect 450 -105 465 -50
rect 480 -60 495 -50
rect 510 -45 555 -35
rect 510 -60 525 -45
rect 540 -60 555 -45
rect 510 -75 555 -60
rect 510 -90 525 -75
rect 510 -100 555 -90
rect 515 -105 555 -100
<< end >>

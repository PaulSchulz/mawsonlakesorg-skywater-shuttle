magic
tech sky130A
timestamp 1598356911
<< metal1 >>
rect 1800 750 1815 855
<< end >>

magic
tech sky130A
timestamp 1598433283
<< metal1 >>
rect 875 850 945 855
rect 870 845 950 850
rect 865 840 955 845
rect 860 835 885 840
rect 935 835 960 840
rect 855 830 880 835
rect 940 830 960 835
rect 855 825 875 830
rect 855 750 870 825
rect 895 820 920 825
rect 890 815 925 820
rect 885 805 930 815
rect 885 770 900 805
rect 915 795 930 805
rect 915 770 930 780
rect 885 760 930 770
rect 890 755 925 760
rect 895 750 920 755
rect 945 750 960 830
rect 855 745 875 750
rect 940 745 960 750
rect 855 740 880 745
rect 935 740 960 745
rect 860 735 885 740
rect 930 735 955 740
rect 865 730 950 735
rect 870 725 945 730
rect 875 720 940 725
<< end >>

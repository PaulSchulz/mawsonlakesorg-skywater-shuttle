magic
tech sky130A
timestamp 1598181805
<< metal1 >>
rect 1135 250 1170 255
rect 1130 245 1170 250
rect 1125 235 1170 245
rect 1125 215 1140 235
rect 1125 210 1160 215
rect 1125 205 1165 210
rect 1130 200 1170 205
rect 1135 195 1170 200
rect 1155 170 1170 195
rect 1125 160 1170 170
rect 1125 155 1165 160
rect 1125 150 1160 155
<< end >>

magic
tech sky130A
timestamp 1598181805
<< metal1 >>
rect 1065 250 1100 255
rect 1065 245 1105 250
rect 1065 235 1110 245
rect 1065 220 1080 235
rect 1095 220 1110 235
rect 1065 210 1110 220
rect 1065 205 1105 210
rect 1065 200 1100 205
rect 1065 185 1095 200
rect 1065 180 1100 185
rect 1065 175 1105 180
rect 1065 165 1110 175
rect 1065 150 1080 165
rect 1095 150 1110 165
<< end >>

magic
tech sky130A
timestamp 1598182001
<< metal1 >>
rect 480 390 525 405
rect 480 375 495 390
rect 510 375 525 390
rect 480 360 525 375
rect 480 315 495 360
rect 510 315 525 360
rect 480 300 525 315
<< end >>

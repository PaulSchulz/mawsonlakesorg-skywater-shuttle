magic
tech sky130A
timestamp 1598363612
<< metal1 >>
rect 1620 450 1650 480
rect 1635 435 1650 450
<< end >>

magic
tech sky130A
timestamp 1598360266
<< metal1 >>
rect -75 795 -15 810
rect -75 765 -15 780
<< end >>

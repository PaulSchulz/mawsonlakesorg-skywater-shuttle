magic
tech sky130A
timestamp 1598177753
<< metal1 >>
rect 320 100 345 105
rect 315 90 345 100
rect 315 75 330 90
rect 300 60 345 75
rect 315 0 330 60
<< end >>

magic
tech sky130A
timestamp 1598181805
<< metal1 >>
rect 1015 250 1040 255
rect 1010 245 1045 250
rect 1005 235 1050 245
rect 1005 185 1020 235
rect 1035 185 1050 235
rect 1005 160 1050 185
rect 1010 155 1050 160
rect 1015 150 1050 155
<< end >>

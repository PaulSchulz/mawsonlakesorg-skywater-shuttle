magic
tech sky130A
timestamp 1598177753
<< metal1 >>
rect 525 75 555 105
rect 525 45 555 60
rect 540 -15 555 45
rect 525 -25 555 -15
rect 525 -30 550 -25
<< end >>

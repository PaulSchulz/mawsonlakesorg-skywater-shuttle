magic
tech sky130A
timestamp 1598356858
<< metal1 >>
rect 1710 825 1740 855
rect 1770 835 1785 855
rect 1765 830 1785 835
rect 1760 825 1785 830
rect 1755 820 1780 825
rect 1755 815 1775 820
rect 1750 810 1770 815
rect 1735 805 1770 810
rect 1730 800 1765 805
rect 1725 795 1760 800
rect 1725 790 1745 795
rect 1720 785 1740 790
rect 1715 780 1740 785
rect 1710 775 1735 780
rect 1710 770 1730 775
rect 1710 750 1725 770
rect 1755 750 1785 780
<< end >>

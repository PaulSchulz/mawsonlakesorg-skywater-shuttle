magic
tech sky130A
timestamp 1598165416
<< metal1 >>
rect 990 70 1025 75
rect 990 65 1030 70
rect 990 55 1035 65
rect 990 0 1005 55
rect 1020 45 1035 55
<< end >>

magic
tech sky130A
timestamp 1598181805
<< metal1 >>
rect 810 240 825 255
rect 810 225 840 240
rect 855 225 870 255
rect 810 210 870 225
rect 810 150 825 210
rect 840 195 870 210
rect 855 150 870 195
<< end >>

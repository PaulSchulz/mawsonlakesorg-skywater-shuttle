magic
tech sky130A
timestamp 1598181805
<< metal1 >>
rect 240 240 285 255
rect 240 210 255 240
rect 240 195 270 210
rect 240 165 255 195
rect 240 150 285 165
<< end >>

magic
tech sky130A
timestamp 1598165416
<< metal1 >>
rect 895 250 920 255
rect 890 245 925 250
rect 885 235 930 245
rect 885 170 900 235
rect 915 170 930 235
rect 885 160 930 170
rect 890 155 925 160
rect 895 150 920 155
<< end >>

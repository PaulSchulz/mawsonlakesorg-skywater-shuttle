magic
tech sky130A
timestamp 1598177753
<< metal1 >>
rect 1380 55 1395 75
rect 1410 55 1425 75
rect 1380 45 1425 55
rect 1385 30 1420 45
rect 1380 20 1425 30
rect 1380 0 1395 20
rect 1410 0 1425 20
<< end >>

magic
tech sky130A
timestamp 1598177753
<< metal1 >>
rect 480 75 510 105
rect 480 45 510 60
rect 495 15 510 45
rect 480 0 510 15
<< end >>

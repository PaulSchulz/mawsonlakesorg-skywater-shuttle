magic
tech sky130A
timestamp 1598165416
<< metal1 >>
rect 370 70 395 75
rect 365 65 400 70
rect 360 55 405 65
rect 360 20 375 55
rect 390 20 405 55
rect 360 10 405 20
rect 365 5 405 10
rect 370 0 405 5
rect 385 -15 405 0
rect 360 -20 405 -15
rect 360 -25 400 -20
rect 360 -30 395 -25
<< end >>

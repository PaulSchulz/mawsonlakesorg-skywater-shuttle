magic
tech sky130A
timestamp 1598359164
<< metal1 >>
rect 1965 845 1990 850
rect 1955 840 1995 845
rect 1950 835 1995 840
rect 2010 835 2025 840
rect 1950 830 2025 835
rect 1950 825 1965 830
rect 1980 825 2025 830
rect 1980 820 2020 825
rect 1985 815 2010 820
<< end >>

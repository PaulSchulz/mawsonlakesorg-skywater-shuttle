magic
tech sky130A
timestamp 1598177753
<< metal1 >>
rect 660 70 690 75
rect 705 70 725 75
rect 660 65 730 70
rect 660 55 735 65
rect 660 0 675 55
rect 690 0 705 55
rect 720 0 735 55
<< end >>

magic
tech sky130A
timestamp 1598362535
<< metal1 >>
rect 2070 820 2085 835
rect 2060 810 2095 820
rect 2045 795 2110 810
rect 2060 785 2095 795
rect 2070 770 2085 785
<< end >>

magic
tech sky130A
timestamp 1598364576
use font_a  font_a_0 lib/font-sky130
timestamp 1598165416
transform 1 0 0 0 1 450
box 0 0 45 75
use font_b  font_b_0 lib/font-sky130
timestamp 1598177753
transform 1 0 0 0 1 450
box 60 0 105 105
use font_c  font_c_0 lib/font-sky130
timestamp 1598177753
transform 1 0 0 0 1 450
box 120 0 165 75
use font_d  font_d_0 lib/font-sky130
timestamp 1598177753
transform 1 0 0 0 1 450
box 180 0 225 105
use font_f  font_f_0 lib/font-sky130
timestamp 1598177753
transform 1 0 0 0 1 450
box 300 0 345 105
use font_e  font_e_0 lib/font-sky130
timestamp 1598165416
transform 1 0 0 0 1 450
box 240 0 285 75
use font_g  font_g_0 lib/font-sky130
timestamp 1598165416
transform 1 0 0 0 1 450
box 360 -30 405 75
use font_h  font_h_0 lib/font-sky130
timestamp 1598177753
transform 1 0 0 0 1 450
box 420 0 465 105
use font_j  font_j_0 lib/font-sky130
timestamp 1598177753
transform 1 0 0 0 1 450
box 525 -30 555 105
use font_i  font_i_0 lib/font-sky130
timestamp 1598177753
transform 1 0 0 0 1 450
box 480 0 510 105
use font_k  font_k_0 lib/font-sky130
timestamp 1598165416
transform 1 0 0 0 1 450
box 570 0 615 105
use font_l  font_l_0 lib/font-sky130
timestamp 1598177753
transform 1 0 0 0 1 450
box 630 0 645 105
use font_m  font_m_0 lib/font-sky130
timestamp 1598177753
transform 1 0 0 0 1 450
box 660 0 735 75
use font_n  font_n_0 lib/font-sky130
timestamp 1598165416
transform 1 0 0 0 1 450
box 750 0 795 75
use font_o  font_o_0 lib/font-sky130
timestamp 1598165416
transform 1 0 0 0 1 450
box 810 0 855 75
use font_p  font_p_0 lib/font-sky130
timestamp 1598177753
transform 1 0 0 0 1 450
box 870 -30 915 75
use font_q  font_q_0 lib/font-sky130
timestamp 1598177753
transform 1 0 0 0 1 450
box 930 -30 975 75
use font_r  font_r_0 lib/font-sky130
timestamp 1598165416
transform 1 0 0 0 1 450
box 990 0 1035 75
use font_s  font_s_0 lib/font-sky130
timestamp 1598165416
transform 1 0 0 0 1 450
box 1050 0 1095 75
use font_t  font_t_0 lib/font-sky130
timestamp 1598177753
transform 1 0 0 0 1 450
box 1110 0 1155 90
use font_u  font_u_0 lib/font-sky130
timestamp 1598177753
transform 1 0 0 0 1 450
box 1170 0 1215 75
use font_v  font_v_0 lib/font-sky130
timestamp 1598177753
transform 1 0 0 0 1 450
box 1230 0 1275 75
use font_w  font_w_0 lib/font-sky130
timestamp 1598166646
transform 1 0 0 0 1 450
box 1290 0 1365 75
use font_2C  font_2C_0 lib/font-sky130
timestamp 1598363612
transform 1 0 0 0 1 0
box 1620 435 1650 480
use font_24  font_24_0 lib/font-sky130
timestamp 1598362656
transform 1 0 0 0 1 0
box 1560 435 1605 540
use font_x  font_x_0 lib/font-sky130
timestamp 1598177753
transform 1 0 0 0 1 450
box 1380 0 1425 75
use font_z  font_z_0 lib/font-sky130
timestamp 1598177753
transform 1 0 0 0 1 450
box 1500 0 1545 75
use font_y  font_y_0 lib/font-sky130
timestamp 1598177753
transform 1 0 0 0 1 450
box 1440 -30 1485 75
use font_01F600  font_01F600_0 lib/font-sky130
timestamp 1598364576
transform 1 0 0 0 1 0
box 1665 450 1770 535
use font_3E  font_3E_0 lib/font-sky130
timestamp 1598360501
transform 1 0 0 0 1 0
box -135 765 -90 840
use font_3C  font_3C_0 lib/font-sky130
timestamp 1598360344
transform 1 0 0 0 1 0
box -195 765 -150 840
use font_B  font_B_0 lib/font-sky130
timestamp 1598181805
transform 1 0 0 0 1 450
box 60 150 105 255
use font_A  font_A_0 lib/font-sky130
timestamp 1598181805
transform 1 0 0 0 1 450
box 0 150 45 255
use font_C  font_C_0 lib/font-sky130
timestamp 1598181805
transform 1 0 0 0 1 450
box 120 150 165 255
use font_0  font_0_0 lib/font-sky130
timestamp 1598182001
transform 1 0 0 0 1 750
box 0 0 45 105
use font_1  font_1_0 lib/font-sky130
timestamp 1598182001
transform 1 0 0 0 1 450
box 60 300 105 405
use font_2  font_2_0 lib/font-sky130
timestamp 1598182001
transform 1 0 0 0 1 450
box 120 300 165 405
use font_3D  font_3D_0 lib/font-sky130
timestamp 1598360266
transform 1 0 0 0 1 15
box -75 765 -15 810
use font_D  font_D_0 lib/font-sky130
timestamp 1598181805
transform 1 0 60 0 1 450
box 120 150 165 255
use font_F  font_F_0 lib/font-sky130
timestamp 1598181805
transform 1 0 0 0 1 450
box 300 150 345 255
use font_E  font_E_0 lib/font-sky130
timestamp 1598181805
transform 1 0 0 0 1 450
box 240 150 285 255
use font_G  font_G_0 lib/font-sky130
timestamp 1598181805
transform 1 0 0 0 1 450
box 360 150 405 255
use font_3  font_3_0 lib/font-sky130
timestamp 1598182472
transform 1 0 0 0 1 450
box 180 300 225 405
use font_5  font_5_0 lib/font-sky130
timestamp 1598182001
transform 1 0 0 0 1 450
box 300 300 345 405
use font_4  font_4_0 lib/font-sky130
timestamp 1598182001
transform 1 0 0 0 1 450
box 240 300 285 405
use font_6  font_6_0 lib/font-sky130
timestamp 1598182001
transform 1 0 0 0 1 450
box 360 300 405 405
use font_3A  font_3A_0 lib/font-sky130
timestamp 1598183786
transform 1 0 0 0 1 0
box 645 750 675 825
use font_2E  font_2E_0 lib/font-sky130
timestamp 1598165416
transform 1 0 -960 0 1 750
box 1560 0 1590 30
use font_H  font_H_0 lib/font-sky130
timestamp 1598181805
transform 1 0 0 0 1 450
box 420 150 465 255
use font_I  font_I_0 lib/font-sky130
timestamp 1598181805
transform 1 0 0 0 1 450
box 480 150 525 255
use font_J  font_J_0 lib/font-sky130
timestamp 1598181805
transform 1 0 0 0 1 450
box 540 150 585 255
use font_K  font_K_0 lib/font-sky130
timestamp 1598181805
transform 1 0 0 0 1 450
box 600 150 645 255
use font_7  font_7_0 lib/font-sky130
timestamp 1598182001
transform 1 0 0 0 1 450
box 420 300 465 405
use font_8  font_8_0 lib/font-sky130
timestamp 1598182001
transform 1 0 0 0 1 450
box 480 300 525 405
use font_9  font_9_0 lib/font-sky130
timestamp 1598182001
transform 1 0 0 0 1 450
box 540 300 585 405
use font_A9  font_A9_0 lib/font-sky130
timestamp 1598185717
transform 1 0 -120 0 1 0
box 855 720 960 855
use font_3B  font_3B_0 lib/font-sky130
timestamp 1598183786
transform 1 0 0 0 1 0
box 690 735 720 825
use font_M  font_M_0 lib/font-sky130
timestamp 1598165416
transform 1 0 0 0 1 450
box 720 150 795 255
use font_L  font_L_0 lib/font-sky130
timestamp 1598165416
transform 1 0 0 0 1 450
box 660 150 705 255
use font_N  font_N_0 lib/font-sky130
timestamp 1598181805
transform 1 0 0 0 1 450
box 810 150 870 255
use font_O  font_O_0 lib/font-sky130
timestamp 1598165416
transform 1 0 0 0 1 450
box 885 150 930 255
use font_40  font_at_0 lib/font-sky130
timestamp 1598185717
transform 1 0 0 0 1 0
box 855 720 960 855
use font_2D  font_2D_0 lib/font-sky130
timestamp 1598355651
transform 1 0 0 0 1 10
box 1065 785 1125 800
use font_21  font_21_0 lib/font-sky130
timestamp 1598361454
transform 1 0 0 0 1 0
box 975 750 1005 855
use font_P  font_P_0 lib/font-sky130
timestamp 1598181805
transform 1 0 0 0 1 450
box 945 150 990 255
use font_Q  font_Q_0 lib/font-sky130
timestamp 1598181805
transform 1 0 0 0 1 450
box 1005 150 1050 255
use font_R  font_R_0 lib/font-sky130
timestamp 1598181805
transform 1 0 0 0 1 450
box 1065 150 1110 255
use font_S  font_S_0 lib/font-sky130
timestamp 1598181805
transform 1 0 0 0 1 450
box 1125 150 1170 255
use font_27  font_27_0 lib/font-sky130
timestamp 1598355651
transform 1 0 0 0 1 0
box 1020 810 1050 855
use font_2B  font_2B_0 lib/font-sky130
timestamp 1598355775
transform 1 0 0 0 1 10
box 1140 770 1185 815
use font_T  font_T_0 lib/font-sky130
timestamp 1598181805
transform 1 0 0 0 1 450
box 1185 150 1230 255
use font_U  font_U_0 lib/font-sky130
timestamp 1598181805
transform 1 0 0 0 1 450
box 1245 150 1290 255
use font_W  font_W_0 lib/font-sky130
timestamp 1598181805
transform 1 0 0 0 1 450
box 1365 150 1440 255
use font_V  font_V_0 lib/font-sky130
timestamp 1598181805
transform 1 0 0 0 1 450
box 1305 150 1350 255
use font_5B  font_5B_0 lib/font-sky130
timestamp 1598356361
transform 1 0 -60 0 1 0
box 1335 750 1380 855
use font_5F  font_5F_0 lib/font-sky130
timestamp 1598356319
transform 1 0 0 0 1 0
box 1200 750 1260 765
use font_5D  font_5D_0 lib/font-sky130
timestamp 1598356419
transform 1 0 -60 0 1 0
box 1395 750 1440 855
use font_X  font_X_0 lib/font-sky130
timestamp 1598181805
transform 1 0 0 0 1 450
box 1455 150 1500 255
use font_Z  font_Z_0 lib/font-sky130
timestamp 1598181805
transform 1 0 0 0 1 450
box 1575 150 1620 255
use font_Y  font_Y_0 lib/font-sky130
timestamp 1598181805
transform 1 0 0 0 1 450
box 1515 150 1560 255
use font_5E  font_5E_0 lib/font-sky130
timestamp 1598356481
transform 1 0 -60 0 1 0
box 1455 825 1500 855
use font_23  font_23_0 lib/font-sky130
timestamp 1598356557
transform 1 0 -60 0 1 0
box 1515 750 1590 855
use font_60  font_60_0 lib/font-sky130
timestamp 1598356612
transform 1 0 -60 0 1 0
box 1605 810 1635 855
use font_2F  font_2F_0 lib/font-sky130
timestamp 1598356782
transform 1 0 -60 0 1 0
box 1650 750 1695 855
use font_3F  font_3F_0 lib/font-sky130
timestamp 1598364457
transform 1 0 0 0 1 0
box 1725 600 1770 705
use font_26  font_26_0 lib/font-sky130
timestamp 1598363904
transform 1 0 0 0 1 0
box 1635 600 1710 705
use font_7D  font_7D_0 lib/font-sky130
timestamp 1598359058
transform 1 0 -60 0 1 0
box 1890 750 1935 855
use font_7B  font_7B_0 lib/font-sky130
timestamp 1598356953
transform 1 0 -60 0 1 0
box 1830 750 1875 855
use font_7C  font_7C_0 lib/font-sky130
timestamp 1598356911
transform 1 0 -60 0 1 0
box 1800 750 1815 855
use font_25  font_25_0 lib/font-sky130
timestamp 1598356858
transform 1 0 -60 0 1 0
box 1710 750 1785 855
use font_2A  font_2A_0 lib/font-sky130
timestamp 1598362535
transform 1 0 -5 0 1 0
box 2045 770 2110 835
use font_22  font_22_0 lib/font-sky130
timestamp 1598359472
transform -1 0 4065 0 1 5
box 2040 790 2085 850
use font_7E  font_7E_0 lib/font-sky130
timestamp 1598359164
transform 1 0 -60 0 1 5
box 1950 815 2025 850
use font_o  font_o_1
timestamp 1598165416
transform 1 0 -750 0 1 960
box 810 0 855 75
use font_F  font_F_1
timestamp 1598181805
transform 1 0 -300 0 1 810
box 300 150 345 255
use font_n  font_n_1
timestamp 1598165416
transform 1 0 -630 0 1 960
box 750 0 795 75
use font_t  font_t_1
timestamp 1598177753
transform 1 0 -930 0 1 960
box 1110 0 1155 90
use font_colon  font_colon_1 lib/font-sky130
timestamp 1598183786
transform 1 0 -405 0 1 210
box 645 750 675 825
use font_s  font_s_1
timestamp 1598165416
transform 1 0 -720 0 1 960
box 1050 0 1095 75
use font_k  font_k_1
timestamp 1598165416
transform 1 0 -180 0 1 960
box 570 0 615 105
use font_1  font_1_1
timestamp 1598182001
transform 1 0 450 0 1 660
box 60 300 105 405
use font_y  font_y_1
timestamp 1598177753
transform 1 0 -990 0 1 960
box 1440 -30 1485 75
use font_3  font_3_1
timestamp 1598182472
transform 1 0 390 0 1 660
box 180 300 225 405
<< properties >>
string FIXED_BBOX -7 -7 52 112
<< end >>

magic
tech sky130A
timestamp 1598177753
<< metal1 >>
rect 420 75 435 105
rect 420 70 455 75
rect 420 65 460 70
rect 420 55 465 65
rect 420 0 435 55
rect 450 0 465 55
<< end >>

magic
tech sky130A
timestamp 1598185717
<< metal1 >>
rect 875 850 945 855
rect 870 845 950 850
rect 865 840 955 845
rect 860 835 885 840
rect 935 835 960 840
rect 855 830 880 835
rect 940 830 960 835
rect 855 825 875 830
rect 855 750 870 825
rect 895 820 920 825
rect 890 815 925 820
rect 885 805 930 815
rect 885 770 900 805
rect 915 770 930 805
rect 945 770 960 830
rect 885 760 960 770
rect 890 755 955 760
rect 895 750 915 755
rect 930 750 950 755
rect 855 745 875 750
rect 855 740 880 745
rect 860 735 885 740
rect 865 730 945 735
rect 870 725 945 730
rect 875 720 945 725
<< end >>

magic
tech sky130A
timestamp 1598355651
<< metal1 >>
rect 1065 785 1125 800
<< end >>

magic
tech sky130A
timestamp 1598165416
<< metal1 >>
rect 570 60 585 105
rect 600 60 615 75
rect 570 50 615 60
rect 570 45 610 50
rect 570 30 600 45
rect 570 25 610 30
rect 570 15 615 25
rect 570 0 585 15
rect 600 0 615 15
<< end >>

magic
tech sky130A
timestamp 1598356953
<< metal1 >>
rect 1855 850 1875 855
rect 1850 845 1875 850
rect 1845 835 1875 845
rect 1845 820 1860 835
rect 1840 810 1860 820
rect 1830 795 1855 810
rect 1840 785 1860 795
rect 1845 770 1860 785
rect 1845 760 1875 770
rect 1850 755 1875 760
rect 1855 750 1875 755
<< end >>

magic
tech sky130A
timestamp 1598181805
<< metal1 >>
rect 1455 230 1470 255
rect 1485 230 1500 255
rect 1455 220 1500 230
rect 1460 210 1495 220
rect 1465 195 1490 210
rect 1460 185 1495 195
rect 1455 175 1500 185
rect 1455 150 1470 175
rect 1485 150 1500 175
<< end >>

magic
tech sky130A
timestamp 1598177753
<< metal1 >>
rect 1230 30 1245 75
rect 1260 30 1275 75
rect 1230 15 1275 30
rect 1235 10 1270 15
rect 1245 0 1260 10
<< end >>

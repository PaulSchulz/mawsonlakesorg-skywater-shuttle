magic
tech sky130A
timestamp 1598181805
<< metal1 >>
rect 1305 205 1320 255
rect 1335 205 1350 255
rect 1305 195 1350 205
rect 1310 180 1345 195
rect 1315 165 1340 180
rect 1320 150 1335 165
<< end >>

magic
tech sky130A
timestamp 1598364457
<< metal1 >>
rect 1735 700 1760 705
rect 1730 695 1765 700
rect 1725 685 1770 695
rect 1725 675 1740 685
rect 1755 665 1770 685
rect 1750 660 1770 665
rect 1740 655 1770 660
rect 1735 650 1765 655
rect 1735 640 1760 650
rect 1730 600 1765 625
<< end >>

magic
tech sky130A
timestamp 1598177753
<< metal1 >>
rect 1440 20 1455 75
rect 1470 20 1485 75
rect 1440 10 1485 20
rect 1445 5 1485 10
rect 1450 0 1485 5
rect 1465 -15 1485 0
rect 1440 -20 1485 -15
rect 1440 -25 1480 -20
rect 1440 -30 1475 -25
<< end >>

magic
tech sky130A
timestamp 1598177753
<< metal1 >>
rect 630 0 645 105
<< end >>

magic
tech sky130A
timestamp 1598181805
<< metal1 >>
rect 1365 205 1380 255
rect 1395 205 1410 255
rect 1425 205 1440 255
rect 1365 195 1440 205
rect 1370 180 1435 195
rect 1375 165 1430 180
rect 1380 150 1395 165
rect 1410 150 1425 165
<< end >>

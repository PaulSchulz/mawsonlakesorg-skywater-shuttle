magic
tech sky130A
timestamp 1598165416
<< metal1 >>
rect 1560 0 1590 30
<< end >>

magic
tech sky130A
timestamp 1598183786
<< metal1 >>
rect 645 795 675 825
rect 645 750 675 780
<< end >>

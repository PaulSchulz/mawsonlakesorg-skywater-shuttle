magic
tech sky130A
timestamp 1598356361
<< metal1 >>
rect 1335 840 1380 855
rect 1335 765 1350 840
rect 1335 750 1380 765
<< end >>

magic
tech sky130A
timestamp 1598355651
<< metal1 >>
rect 1020 825 1050 855
rect 1035 810 1050 825
<< end >>

magic
tech sky130A
timestamp 1598165416
<< metal1 >>
rect 820 70 845 75
rect 815 65 850 70
rect 810 55 855 65
rect 810 20 825 55
rect 840 20 855 55
rect 810 10 855 20
rect 815 5 850 10
rect 820 0 845 5
<< end >>

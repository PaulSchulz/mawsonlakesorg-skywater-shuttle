magic
tech sky130A
timestamp 1598356419
<< metal1 >>
rect 1395 840 1440 855
rect 1425 765 1440 840
rect 1395 750 1440 765
<< end >>

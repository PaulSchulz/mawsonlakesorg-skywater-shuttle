magic
tech sky130A
timestamp 1598181805
<< metal1 >>
rect 1515 220 1530 255
rect 1545 220 1560 255
rect 1515 210 1560 220
rect 1520 200 1555 210
rect 1525 190 1550 200
rect 1530 150 1545 190
<< end >>

magic
tech sky130A
timestamp 1598181805
<< metal1 >>
rect 480 240 525 255
rect 495 165 510 240
rect 480 150 525 165
<< end >>

magic
tech sky130A
timestamp 1598185717
<< metal1 >>
rect 755 850 820 855
rect 750 845 825 850
rect 745 840 830 845
rect 740 835 765 840
rect 810 835 835 840
rect 735 830 760 835
rect 815 830 840 835
rect 735 825 755 830
rect 820 825 840 830
rect 735 750 750 825
rect 775 820 800 825
rect 770 815 805 820
rect 765 805 810 815
rect 765 770 780 805
rect 795 795 810 805
rect 795 770 810 780
rect 765 760 810 770
rect 770 755 805 760
rect 775 750 800 755
rect 825 750 840 825
rect 735 745 755 750
rect 820 745 840 750
rect 735 740 760 745
rect 815 740 840 745
rect 740 735 765 740
rect 810 735 835 740
rect 745 730 830 735
rect 750 725 825 730
rect 755 720 820 725
<< end >>

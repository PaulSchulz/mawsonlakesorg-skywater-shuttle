magic
tech sky130A
timestamp 1598177753
<< metal1 >>
rect 1125 75 1140 90
rect 1110 60 1155 75
rect 1125 0 1140 60
<< end >>

magic
tech sky130A
timestamp 1598356612
<< metal1 >>
rect 1605 825 1635 855
rect 1605 810 1620 825
<< end >>
